module hello_world

pub fn say() string {
	return 'Hello, world!'
}
