module helloworld

pub fn say() string {
	return 'Hello, world!'
}
