module main

fn test_hello() {
	assert say() == 'Hello, world!'
}
