module hello_world

pub fn say() string {
  return "Goodbye, world!"
}
