module main

fn say() string {
	return 'Goodbye, world!'
}
