module hello_world_mismatched

pub fn say() string {
	return 'Hello, world!'
}
