module helloworld

pub fn say() string {
	return 'Goodbye, world!'
}
