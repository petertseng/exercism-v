module hello-world

pub fn say() string {
  return "Hello, world!"
}
