module main

fn leap(year int) bool {
  panic("determine whether the year is a leap year")
}
