module main

fn say() string {
	return 'Hello, world!'
}
