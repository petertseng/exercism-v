module hello-world

pub fn say() string {
  return "Goodbye, world!"
}
